Embedded_Multiplier_16_inst : Embedded_Multiplier_16 PORT MAP (
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		result	 => result_sig
	);
